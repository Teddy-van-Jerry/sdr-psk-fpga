module Not_Gate (
  input  i,
  output o
);
  assign o = ~i; 
endmodule
